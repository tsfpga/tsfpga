// -------------------------------------------------------------------------------------------------
// Copyright (c) Lukas Vik. All rights reserved.
//
// This file is part of the tsfpga project, a project platform for modern FPGA development.
// https://tsfpga.com
// https://github.com/tsfpga/tsfpga
// -------------------------------------------------------------------------------------------------

package artyz7_top_systemverilog_pkg;

  localparam int num_leds = 4;

endpackage : artyz7_top_systemverilog_pkg
